module InstMem(PC, instruction);
input [31:0] PC;
output [31:0] instruction;
reg[31:0] memory[0:19];
initial
    begin
        memory[0] <= 32'b00111001100100000000001100010011;
		memory[1] <= 32'b00000000011000000010001000100011;
		memory[2] <= 32'b00000000010000000000001010000011;
		memory[3] <= 32'b00000000010100000010000000100011;
		memory[4] <= 32'b00000010000000110000000001100011;
		memory[5] <= 32'b00000000000000000010111000000011;
		memory[6] <= 32'b00000001110000101001110001100011;
		memory[7] <= 32'b00000001110000101000001110110011;
		memory[8] <= 32'b00000001110000111111001100110011;
		memory[9] <= 32'b00000000000000111111001100010011;
		memory[10] <= 32'b01000000000000110000001010110011;
		memory[11] <= 32'b00000000011000101101010001100011;
		memory[12] <= 32'b00000000000000000000001110110011;
		memory[13] <= 32'b00000000110000000000000011101111;
		memory[14] <= 32'b00000001010000000000000011101111;
		memory[15] <= 32'b00000000000000000000111000110011;
		memory[16] <= 32'b00000000011111100110111000110011;
		memory[17] <= 32'b00000000000000001000000001100111;
		memory[18] <= 32'b00000100100000000000001100010011;
		memory[19] <= 32'b00001010110000000000001010010011;
    end
assign instruction=memory[PC>>2];
endmodule
